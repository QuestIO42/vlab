module top(input [3:0] SW, output [3:0] LEDR);
	assign LEDR = SW;
endmodule 
